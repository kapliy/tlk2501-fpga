library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity disparity_lookup is
	port
	(
		clk_in : in STD_LOGIC;
		data_in : in STD_LOGIC_VECTOR(7 downto 0);
		dispflip_out : out STD_LOGIC
	);
end disparity_lookup;

architecture structure of disparity_lookup is

type TYPE_DISPFLIP_LUP is array (0 to 255) of STD_LOGIC;
-- 02/19/2011 - changed lup from "signal" to "constant"
constant DISPFLIP_LUP : TYPE_DISPFLIP_LUP:=
          (
          '0', -- "00000000"
          '0', -- "00000001"
          '0', -- "00000010"
          '1', -- "00000011"
          '0', -- "00000100"
          '1', -- "00000101"
          '1', -- "00000110"
          '1', -- "00000111"
          '0', -- "00001000"
          '1', -- "00001001"
          '1', -- "00001010"
          '1', -- "00001011"
          '1', -- "00001100"
          '1', -- "00001101"
          '1', -- "00001110"
          '0', -- "00001111"
          '0', -- "00010000"
          '1', -- "00010001"
          '1', -- "00010010"
          '1', -- "00010011"
          '1', -- "00010100"
          '1', -- "00010101"
          '1', -- "00010110"
          '0', -- "00010111"
          '0', -- "00011000"
          '1', -- "00011001"
          '1', -- "00011010"
          '0', -- "00011011"
          '1', -- "00011100"
          '0', -- "00011101"
          '0', -- "00011110"
          '0', -- "00011111"
          '1', -- "00100000"
          '1', -- "00100001"
          '1', -- "00100010"
          '0', -- "00100011"
          '1', -- "00100100"
          '0', -- "00100101"
          '0', -- "00100110"
          '0', -- "00100111"
          '1', -- "00101000"
          '0', -- "00101001"
          '0', -- "00101010"
          '0', -- "00101011"
          '0', -- "00101100"
          '0', -- "00101101"
          '0', -- "00101110"
          '1', -- "00101111"
          '1', -- "00110000"
          '0', -- "00110001"
          '0', -- "00110010"
          '0', -- "00110011"
          '0', -- "00110100"
          '0', -- "00110101"
          '0', -- "00110110"
          '1', -- "00110111"
          '1', -- "00111000"
          '0', -- "00111001"
          '0', -- "00111010"
          '1', -- "00111011"
          '0', -- "00111100"
          '1', -- "00111101"
          '1', -- "00111110"
          '1', -- "00111111"
          '1', -- "01000000"
          '1', -- "01000001"
          '1', -- "01000010"
          '0', -- "01000011"
          '1', -- "01000100"
          '0', -- "01000101"
          '0', -- "01000110"
          '0', -- "01000111"
          '1', -- "01001000"
          '0', -- "01001001"
          '0', -- "01001010"
          '0', -- "01001011"
          '0', -- "01001100"
          '0', -- "01001101"
          '0', -- "01001110"
          '1', -- "01001111"
          '1', -- "01010000"
          '0', -- "01010001"
          '0', -- "01010010"
          '0', -- "01010011"
          '0', -- "01010100"
          '0', -- "01010101"
          '0', -- "01010110"
          '1', -- "01010111"
          '1', -- "01011000"
          '0', -- "01011001"
          '0', -- "01011010"
          '1', -- "01011011"
          '0', -- "01011100"
          '1', -- "01011101"
          '1', -- "01011110"
          '1', -- "01011111"
          '1', -- "01100000"
          '1', -- "01100001"
          '1', -- "01100010"
          '0', -- "01100011"
          '1', -- "01100100"
          '0', -- "01100101"
          '0', -- "01100110"
          '0', -- "01100111"
          '1', -- "01101000"
          '0', -- "01101001"
          '0', -- "01101010"
          '0', -- "01101011"
          '0', -- "01101100"
          '0', -- "01101101"
          '0', -- "01101110"
          '1', -- "01101111"
          '1', -- "01110000"
          '0', -- "01110001"
          '0', -- "01110010"
          '0', -- "01110011"
          '0', -- "01110100"
          '0', -- "01110101"
          '0', -- "01110110"
          '1', -- "01110111"
          '1', -- "01111000"
          '0', -- "01111001"
          '0', -- "01111010"
          '1', -- "01111011"
          '0', -- "01111100"
          '1', -- "01111101"
          '1', -- "01111110"
          '1', -- "01111111"
          '0', -- "10000000"
          '0', -- "10000001"
          '0', -- "10000010"
          '1', -- "10000011"
          '0', -- "10000100"
          '1', -- "10000101"
          '1', -- "10000110"
          '1', -- "10000111"
          '0', -- "10001000"
          '1', -- "10001001"
          '1', -- "10001010"
          '1', -- "10001011"
          '1', -- "10001100"
          '1', -- "10001101"
          '1', -- "10001110"
          '0', -- "10001111"
          '0', -- "10010000"
          '1', -- "10010001"
          '1', -- "10010010"
          '1', -- "10010011"
          '1', -- "10010100"
          '1', -- "10010101"
          '1', -- "10010110"
          '0', -- "10010111"
          '0', -- "10011000"
          '1', -- "10011001"
          '1', -- "10011010"
          '0', -- "10011011"
          '1', -- "10011100"
          '0', -- "10011101"
          '0', -- "10011110"
          '0', -- "10011111"
          '1', -- "10100000"
          '1', -- "10100001"
          '1', -- "10100010"
          '0', -- "10100011"
          '1', -- "10100100"
          '0', -- "10100101"
          '0', -- "10100110"
          '0', -- "10100111"
          '1', -- "10101000"
          '0', -- "10101001"
          '0', -- "10101010"
          '0', -- "10101011"
          '0', -- "10101100"
          '0', -- "10101101"
          '0', -- "10101110"
          '1', -- "10101111"
          '1', -- "10110000"
          '0', -- "10110001"
          '0', -- "10110010"
          '0', -- "10110011"
          '0', -- "10110100"
          '0', -- "10110101"
          '0', -- "10110110"
          '1', -- "10110111"
          '1', -- "10111000"
          '0', -- "10111001"
          '0', -- "10111010"
          '1', -- "10111011"
          '0', -- "10111100"
          '1', -- "10111101"
          '1', -- "10111110"
          '1', -- "10111111"
          '1', -- "11000000"
          '1', -- "11000001"
          '1', -- "11000010"
          '0', -- "11000011"
          '1', -- "11000100"
          '0', -- "11000101"
          '0', -- "11000110"
          '0', -- "11000111"
          '1', -- "11001000"
          '0', -- "11001001"
          '0', -- "11001010"
          '0', -- "11001011"
          '0', -- "11001100"
          '0', -- "11001101"
          '0', -- "11001110"
          '1', -- "11001111"
          '1', -- "11010000"
          '0', -- "11010001"
          '0', -- "11010010"
          '0', -- "11010011"
          '0', -- "11010100"
          '0', -- "11010101"
          '0', -- "11010110"
          '1', -- "11010111"
          '1', -- "11011000"
          '0', -- "11011001"
          '0', -- "11011010"
          '1', -- "11011011"
          '0', -- "11011100"
          '1', -- "11011101"
          '1', -- "11011110"
          '1', -- "11011111"
          '0', -- "11100000"
          '0', -- "11100001"
          '0', -- "11100010"
          '1', -- "11100011"
          '0', -- "11100100"
          '1', -- "11100101"
          '1', -- "11100110"
          '1', -- "11100111"
          '0', -- "11101000"
          '1', -- "11101001"
          '1', -- "11101010"
          '1', -- "11101011"
          '1', -- "11101100"
          '1', -- "11101101"
          '1', -- "11101110"
          '0', -- "11101111"
          '0', -- "11110000"
          '1', -- "11110001"
          '1', -- "11110010"
          '1', -- "11110011"
          '1', -- "11110100"
          '1', -- "11110101"
          '1', -- "11110110"
          '0', -- "11110111"
          '0', -- "11111000"
          '1', -- "11111001"
          '1', -- "11111010"
          '0', -- "11111011"
          '1', -- "11111100"
          '0', -- "11111101"
          '0', -- "11111110"
          '0'  -- "11111111"
);

signal dispflip : STD_LOGIC;
begin
  dispflip_out <= dispflip;

  -- the following LUT might be synthesized into a ROM memory (altsyncram)
  process (clk_in)
  begin
    if (clk_in='1' and clk_in'event)
    then
      dispflip <= DISPFLIP_LUP(conv_integer(data_in));
    end if;
  end process;
end structure;
